--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   11:50:54 05/11/2012
-- Design Name:   
-- Module Name:   C:/Xilinx/dige1/avr_keypad/tb_decoder_columns.vhd
-- Project Name:  avr_keypad
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: decoder_columns
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_decoder_columns IS
END tb_decoder_columns;
 
ARCHITECTURE behavior OF tb_decoder_columns IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT decoder_columns
    PORT(
         dec_in : IN  std_logic_vector(1 downto 0);
         dec_out : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal dec_in : std_logic_vector(1 downto 0) := (others => '0');

 	--Outputs
   signal dec_out : std_logic_vector(3 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: decoder_columns PORT MAP (
          dec_in => dec_in,
          dec_out => dec_out
        );



   -- Stimulus process
   stim_proc: process
   begin		
    
	 wait for 100 ns;
		dec_in <= "00";		-- dec_out must be 0001
	 wait for 100 ns;
		dec_in <= "01"; 		-- dec_out must be 0010
	 wait for 100 ns;
		dec_in <= "10"; 		-- dec_out must be 0100
	 wait for 100 ns;
		dec_in <= "11"; 		-- dec_out must be 1000
	 
	 
      wait;
   end process;

END;
