`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:53:40 05/25/2012 
// Design Name: 
// Module Name:    key_press 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module key_press(
    input [3:0] in_keypad,
    input en_cnt,
    input rst_cnt,
    input [3:0] in_col,
    output [4:0] btn_press
    );


endmodule
